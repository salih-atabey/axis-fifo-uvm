package axis_if_pkg;
    parameter integer DATA_WIDTH = 64;
    parameter integer ID_WIDTH = 8;
    parameter integer DEST_WIDTH = 8;
    parameter integer USER_WIDTH = 8;
endpackage
